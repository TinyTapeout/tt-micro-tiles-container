// Just a stub to make tests happy

`default_nettype none

module tt_um_watbulb_sync_fifo (
    input  wire [7:0] ui_in,   // Dedicated inputs
    output wire [7:0] uo_out,  // Dedicated outputs
    input  wire       clk,     // clock
    input  wire       rst_n    // reset_n - low to reset
);

endmodule
